module PhaseCounter(
    
);
// 在此次设计中，2pai分解为256个点
endmodule   // PhaseCounter